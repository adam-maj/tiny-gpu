`default_nettype none
`timescale 1ns/1ns

// ARITHMETIC-LOGIC UNIT
module alu (
    // Control
    input wire clk,
    input wire reset,
)

endmodule