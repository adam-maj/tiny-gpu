`default_nettype none
`timescale 1ns/1ns

// L1 CACHE
module cache (
    // Control
    input wire clk,
    input wire reset,
)

endmodule