`default_nettype none
`timescale 1ns/1ns

// DISPATCHER
module dispatcher (
    // Control
    input wire clk,
    input wire reset,
);

endmodule