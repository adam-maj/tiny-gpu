`default_nettype none
`timescale 1ns/1ns

// ISSUER
module issuer (
    // Control
    input wire clk,
    input wire reset,
)

endmodule