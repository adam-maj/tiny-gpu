`default_nettype none
`timescale 1ns/1ns

// WARP SCHEDULER
module warps (
    // Control
    input wire clk,
    input wire reset,
)
    // DAG

    // Reservation Station / Scoreboard
endmodule