`default_nettype none
`timescale 1ns/1ns

// DECODER
module decoder (
    // Control
    input wire clk,
    input wire reset,
)

endmodule