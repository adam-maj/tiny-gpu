`default_nettype none
`timescale 1ns/1ns

// REGISTER FILE
module registers (
    // Control
    input wire clk,
    input wire reset,
)

endmodule