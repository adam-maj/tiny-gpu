`default_nettype none
`timescale 1ns/1ns

// STREAMING MULTI-PROCESSOR
module sm (
    // Control
    input wire clk,
    input wire reset,

    // Input
    input wire program_counter,
    input wire thread_count,
);
    // === MEMORY === ///

    // Register File

    // L1 Cache
    
    // === LOGIC === //

    // Fetcher

    // Decoder

    // Warp Scheduler

    // Issuer
endmodule

