`default_nettype none
`timescale 1ns/1ns

// FETCHER
module fetcher (
    // Control
    input wire clk,
    input wire reset,
)

endmodule